
--17030140002 5.11 test4 data-conversion

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity lut is

end lut;

architecture Behavioral of lut is

begin


end Behavioral;

